`include "uvm_macros.svh"
package tb_pkg;
  import uvm_pkg::*;
  `include "transaction.sv"
  `include "sequence.sv"
  `include "sequencer.sv"
  `include "driver.sv"
  `include 'monitor.sv"
  `include "agent.sv"
  `include "predictor.sv"
  `include "comparator.sv"
  `include "scoreboard.sv"
  `include "environment.sv"
  `include "base_test.sv"
endpackage
